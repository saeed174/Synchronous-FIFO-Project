package shared_pkg;

    logic test_finished = 0;
    int correct_count = 0, error_count = 0;
    event driver_finished;

endpackage